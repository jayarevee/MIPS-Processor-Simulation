
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DFlip is
port(D: in STD_LOGIC;
	Clk: in std_logic;
	Reset:in STD_LOGIC;
	Q:out STD_LOGIC
	);
end DFlip;

architecture Behavioral of DFlip is

begin
	process (clk) is
	begin
	if rising_edge(clk) then
		if(reset = '1') then
			Q <= '0';
		
		else
			Q <= D;
		end if;
	end if;
	end process;
end Behavioral;

